RC Circuit
.include vin_piecewise.spice.in
r1 1 2 1MEG
c1 2 0 1uF
.ic V(1)=0 V(2)=0
.tran .001s 5s
.end

